rom_256_x8_lab8_inst : rom_256_x8_lab8 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
