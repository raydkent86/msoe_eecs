rom_64k_x16_v2_inst : rom_64k_x16_v2 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
