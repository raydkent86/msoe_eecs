rom_64k_x16_inst : rom_64k_x16 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
